/********************************************************************
*																	*
*	Boundary_Scan_Cell:												*
*																	*
*	data_in:  values that come from on-chip logic and goes to chip 	*
*	data_out: values that is goes to core							*
*	scan_in: values from previous cell or TDI  						*
*	scan_out: values for next cell or TDO							*
*	ClockDR: Test Clock Generated by Tap Controller					*
*	ShiftDR, UpdateDR: TAP States									*
*	mode: EXTEST or INTEST											*
*																	*
*																	*
********************************************************************/

`timescale 1ns/100ps

module Boundary_Scan_Cell(data_in, data_out, scan_in, scan_out, ClockDR, ShiftDR, UpdateDR, mode);
parameter SIZE = 4;
	
//input
input [SIZE-1:0] data_in;
input scan_in;

//output
output [SIZE-1:0] data_out;
output reg scan_out;

//control signal
input ClockDR;
input ShiftDR;
input UpdateDR;
input mode;


reg	[SIZE-1 : 0] BSC_Scan_Register, BSC_Output_Register;

always @ (posedge ClockDR) begin
	BSC_Scan_Register <= ShiftDR ? {scan_in, BSC_Scan_Register[SIZE-1: 1]} : data_in;
end

always @ (posedge UpdateDR) begin
	BSC_Output_Register <= BSC_Scan_Register;
end

assign scan_out = BSC_Scan_Register [0];
assign data_out = mode ? BSC_Output_Register : data_in;
	

endmodule